module main_mem_controller

	(
		inout			[31:0]			DATA_DQ,
		output			[19:0]			SRAM_ADDR,
		output						SRAM_CE_N, SRAM_OE_N, SRAM_WE_N, SRAM_UB_N, SRAM_LB_N,
		input						clk
	);

	

endmodule
